
typedef enum bit {
    OBI_COV_ENABLE , 
    OBI_COV_DISABLE
} obi_cov_enable_enum;

typedef enum int {
    OBI_RST_STATE_PRE_RESET ,
    OBI_RST_STATE_IN_RESET  ,
    OBI_RST_STATE_POST_RESET
} obi_reset_state_enum;
