
`define RISCV_FORMAL
`define RISCV_FORMAL_NRET 1
`define RISCV_FORMAL_XLEN 32
`define RISCV_FORMAL_ILEN 32
`define RISCV_FORMAL_CSR_MARCHID
`define RISCV_FORMAL_CSR_MCAUSE
`define RISCV_FORMAL_CSR_MEPC
`define RISCV_FORMAL_CSR_MHARTID
`define RISCV_FORMAL_CSR_MIE
`define RISCV_FORMAL_CSR_MIMPID
`define RISCV_FORMAL_CSR_MISA
`define RISCV_FORMAL_CSR_MSTATUS
`define RISCV_FORMAL_CSR_MTVEC
`define RISCV_FORMAL_CSR_MVENDORID
`include "rvfi_macros.vh"