typedef enum bit {
    RVVI_COV_ENABLE , 
    RVVI_COV_DISABLE
} rvvi_cov_enable_enum;

typedef enum bit {
    RVVI_LOGGING_ENABLE , 
    RVVI_LOGGING_DISABLE
} rvvi_logging_enable_enum;
