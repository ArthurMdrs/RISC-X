module rvfi import core_pkg::*; (
    input  logic clk_i,
    input  logic rst_n_i,
    
    // Input from IF stage
    input  logic         valid_if,
    input  logic         stall_if,
    input  logic [31:0]  pc_if,
    input  next_pc_mux_t next_pc_mux,
    
    // Input from ID stage
    input  logic          valid_id,
    input  logic          stall_id,
    input  logic          flush_id,
    input  logic          trap_id,
    input  logic [31:0]   instr_id,
    input  logic          illegal_instr_id,
    input  alu_source_1_t alu_source_1_id,
    input  alu_source_2_t alu_source_2_id,
    input  logic [ 4:0]   rs1_addr_id,
    input  logic [ 4:0]   rs2_addr_id,
    // input  logic [ 4:0]   rs3_addr_id,
    input  reg_bank_mux_t rs1_src_bank_id,
    input  reg_bank_mux_t rs2_src_bank_id,
    input  reg_bank_mux_t rs3_src_bank_id,
    input  logic [31:0]   rs1_or_fwd_id,
    input  logic [31:0]   rs2_or_fwd_id,
    input  logic [31:0]   pc_id,
    input  pc_source_t    pc_source_id,
    input  logic [31:0]   jump_target_id,
    input  logic          mem_wen_id,
    
    // Input from EX stage
    input  logic           valid_ex,
    input  logic           stall_ex,
    input  logic           flush_ex,
    input  logic           trap_ex,
    input  logic [31:0]    branch_target_ex,
    input  logic           branch_decision_ex,
    input  logic [31:0]    csr_wdata_ex,
    input  logic [31:0]    csr_rdata_ex,
    input  csr_operation_t csr_op_ex,
    
    // Input from MEM stage
    input  logic        valid_mem,
    input  logic        stall_mem,
    input  logic        flush_mem,
    input  logic [31:0] dmem_wdata_o,
    input  logic [31:0] dmem_addr_o,
    input  logic        dmem_wen_o,
    input  logic [ 3:0] dmem_ben_o,
    
    // Input from WB stage
    input  logic          flush_wb,
    input  logic [ 4:0]   rd_addr_wb,
    input  reg_bank_mux_t rd_dst_bank_wb,
    input  logic          reg_wen_wb,
    input  logic [31:0]   reg_wdata_wb,
    input  logic [31:0]   mem_rdata_wb,
    
    input  logic [31:0] misa,
    
    `RVFI_OUTPUTS
);

logic        intr_if;

// logic        rvfi_valid_id;
logic        intr_id;

// logic        rvfi_valid_ex;
logic [31:0] instr_ex;
logic        rvfi_trap_ex;
logic        intr_ex;
logic [ 4:0] rs1_addr_ex, rs2_addr_ex;
logic [31:0] rs1_rdata_ex, rs2_rdata_ex;
logic [31:0] pc_ex, pc_n_ex;

// logic        rvfi_valid_mem;
logic [31:0] instr_mem;
logic        trap_mem;
logic        intr_mem;
logic [ 4:0] rs1_addr_mem, rs2_addr_mem;
logic [31:0] rs1_rdata_mem, rs2_rdata_mem;
logic [31:0] pc_mem, pc_n_mem;
logic [31:0] csr_wdata_mem, csr_rdata_mem;
logic        csr_wen_mem;

logic        rvfi_valid_wb;
logic [63:0] order_wb;
logic [31:0] instr_wb;
logic        trap_wb;
logic        intr_wb;
logic [ 4:0] rs1_addr_wb, rs2_addr_wb;
logic [31:0] rs1_rdata_wb, rs2_rdata_wb;
logic [31:0] pc_wb, pc_n_wb;
logic [31:0] mem_addr_wb;
logic [ 3:0] mem_wmask_wb, mem_rmask_wb;
logic [31:0] mem_wdata_wb;//, mem_rdata_wb;
logic [31:0] csr_wdata_wb, csr_rdata_wb;
logic        csr_wen_wb;

`default_nettype none

///////////////////////////////////////////////////////////////////////////////
//////////////////////        INSTRUCTION FETCH         ///////////////////////
///////////////////////////////////////////////////////////////////////////////

// Pipeline registers ->IF
always_ff @(posedge clk_i, negedge rst_n_i) begin
    if (!rst_n_i) begin
        intr_if <= '0;
    end else begin
        if (!stall_if) begin
            intr_if <= (next_pc_mux == NPC_EXCEPTION);
        end
    end
end

///////////////////////////////////////////////////////////////////////////////
//////////////////////        INSTRUCTION DECODE        ///////////////////////
///////////////////////////////////////////////////////////////////////////////

// Pipeline registers IF->ID
always_ff @(posedge clk_i, negedge rst_n_i) begin
    if (!rst_n_i) begin
        // rvfi_valid_id <= '0;
        intr_id <= '0;
    end else begin
        if (!stall_id) begin
            // Insert bubble if flushing is needed
            if (flush_id) begin
                // rvfi_valid_id <= 1'b0;
                intr_id <= '0;
            end
            else begin
                // rvfi_valid_id <= 1'b1;
                intr_id <= intr_if;
            end
        end
    end
end

///////////////////////////////////////////////////////////////////////////////
/////////////////////////           EXECUTE           /////////////////////////
///////////////////////////////////////////////////////////////////////////////

// Pipeline registers ID->EX
always_ff @(posedge clk_i, negedge rst_n_i) begin
    if (!rst_n_i) begin
        // rvfi_valid_ex <= '0;
        instr_ex      <= '0;
        rvfi_trap_ex  <= '0;
        intr_ex       <= '0;
        rs1_addr_ex   <= '0;
        rs2_addr_ex   <= '0;
        rs1_rdata_ex  <= '0;
        rs2_rdata_ex  <= '0;
        pc_ex         <= '0;
        pc_n_ex       <= '0;
    end else begin
        if (!stall_ex) begin
            // instr_ex     <= instr_id;
            instr_ex     <= (instr_id[1:0] == 2'b11) ? (instr_id) : ({16'b0, instr_id[15:0]});
            rvfi_trap_ex <= trap_id && !stall_id && !branch_decision_ex;
            intr_ex      <= intr_id;
            // TODO: use signal rs1_is_used from decoder (when it's implemented)
            if ((rs1_src_bank_id == X_REG) && ((alu_source_1_id == ALU_SCR1_RS1) || (pc_source_id == PC_JALR))) begin
                rs1_addr_ex  <= rs1_addr_id;
                rs1_rdata_ex <= rs1_or_fwd_id;
            end else begin
                rs1_addr_ex  <= '0;
                rs1_rdata_ex <= '0;
            end
            if ((rs2_src_bank_id == X_REG) && ((alu_source_2_id == ALU_SCR2_RS2) || mem_wen_id)) begin
                rs2_addr_ex  <= rs2_addr_id;
                rs2_rdata_ex <= rs2_or_fwd_id;
            end else begin
                rs2_addr_ex  <= '0;
                rs2_rdata_ex <= '0;
            end
            pc_ex        <= pc_id;
            // pc_n_ex <= (pc_source_id inside {PC_JAL, PC_JALR}) ? (jump_target_id) : (pc_if);
            // Insert bubble if flushing is needed
            if (flush_ex) begin
                pc_n_ex       <= '0;
            end
            else begin
                pc_n_ex <= (pc_source_id inside {PC_JAL, PC_JALR}) ? (jump_target_id) : (pc_if);
            end
        end
    end
end

///////////////////////////////////////////////////////////////////////////////
///////////////////////          MEMORY ACCESS          ///////////////////////
///////////////////////////////////////////////////////////////////////////////

// Pipeline registers EX->MEM
always_ff @(posedge clk_i, negedge rst_n_i) begin
    if (!rst_n_i) begin
        // rvfi_valid_mem <= '0;
        instr_mem      <= '0;
        trap_mem       <= '0;
        intr_mem       <= '0;
        rs1_addr_mem   <= '0;
        rs2_addr_mem   <= '0;
        rs1_rdata_mem  <= '0;
        rs2_rdata_mem  <= '0;
        pc_mem         <= '0;
        pc_n_mem       <= '0;
        csr_wdata_mem  <= '0;
        csr_rdata_mem  <= '0;
        csr_wen_mem    <= '0;
    end else begin
        if (!stall_mem) begin
            instr_mem      <= instr_ex;
            trap_mem <= rvfi_trap_ex || (trap_ex && !stall_ex);
            intr_mem <= intr_ex;
            rs1_addr_mem   <= rs1_addr_ex;
            rs2_addr_mem   <= rs2_addr_ex;
            rs1_rdata_mem  <= rs1_rdata_ex;
            rs2_rdata_mem  <= rs2_rdata_ex;
            pc_mem   <= pc_ex;
            // pc_n_mem <= (branch_decision_ex) ? (branch_target_ex) : (pc_n_ex);
            // Insert bubble if flushing is needed
            if (flush_mem) begin
                pc_n_mem       <= '0;    
                csr_wdata_mem  <= '0;
                csr_rdata_mem  <= '0;
                csr_wen_mem    <= '0;
            end
            else begin
                pc_n_mem       <= (branch_decision_ex) ? (branch_target_ex) : (pc_n_ex);
                csr_wdata_mem  <= csr_wdata_ex;
                csr_rdata_mem  <= csr_rdata_ex;
                csr_wen_mem    <= (csr_op_ex != CSR_READ);
            end
        end
    end
end

///////////////////////////////////////////////////////////////////////////////
////////////////////////          WRITE BACK          /////////////////////////
///////////////////////////////////////////////////////////////////////////////

// Pipeline registers EX->MEM
always_ff @(posedge clk_i, negedge rst_n_i) begin
    if (!rst_n_i) begin
        rvfi_valid_wb <= '0;
        order_wb      <= '0;
        instr_wb      <= '0;
        trap_wb       <= '0;
        intr_wb       <= '0;
        rs1_addr_wb   <= '0;
        rs2_addr_wb   <= '0;
        rs1_rdata_wb  <= '0;
        rs2_rdata_wb  <= '0;
        pc_wb         <= '0;
        pc_n_wb       <= '0;
        mem_addr_wb   <= '0;
        mem_rmask_wb  <= '0;
        mem_wmask_wb  <= '0;
        mem_wdata_wb  <= '0;
        csr_wdata_wb  <= '0;
        csr_rdata_wb  <= '0;
        csr_wen_wb    <= '0;
    end else begin
        order_wb <= order_wb + {63'b0, rvfi_valid};
        instr_wb      <= instr_mem;
        trap_wb  <= trap_mem;
        intr_wb  <= intr_mem;
        rs1_addr_wb   <= rs1_addr_mem;
        rs2_addr_wb   <= rs2_addr_mem;
        rs1_rdata_wb  <= rs1_rdata_mem;
        rs2_rdata_wb  <= rs2_rdata_mem;
        pc_wb    <= pc_mem;
        // pc_n_wb  <= pc_n_mem;
        // Insert bubble if flushing is needed
        if (flush_wb) begin
            rvfi_valid_wb <= '0;
            pc_n_wb       <= '0;
            mem_addr_wb   <= '0;
            mem_rmask_wb  <= '0;
            mem_wmask_wb  <= '0;
            mem_wdata_wb  <= '0;
            csr_wdata_wb  <= '0;
            csr_rdata_wb  <= '0;
            csr_wen_wb    <= '0;
        end
        else begin
            // rvfi_valid_wb <= rvfi_valid_mem;
            rvfi_valid_wb <= valid_mem;
            pc_n_wb       <= pc_n_mem;
            mem_addr_wb   <= dmem_addr_o;
            mem_rmask_wb  <= dmem_ben_o;
            mem_wmask_wb  <= (dmem_wen_o) ? (dmem_ben_o) : ('0);
            mem_wdata_wb  <= dmem_wdata_o;
            csr_wdata_wb  <= csr_wdata_mem;
            csr_rdata_wb  <= csr_rdata_mem;
            csr_wen_wb    <= csr_wen_mem;
        end
    end
end

///////////////////////////////////////////////////////////////////////////////
////////////////////////             RVFI             /////////////////////////
///////////////////////////////////////////////////////////////////////////////

// Instruction Metadata
assign rvfi_valid = rvfi_valid_wb || trap_wb;
assign rvfi_order = order_wb;
assign rvfi_insn = instr_wb;
assign rvfi_trap = trap_wb;
assign rvfi_halt = 1'b0;
assign rvfi_intr = intr_wb;
assign rvfi_mode = 2'b11;
assign rvfi_ixl  = 2'b01;

// Integer Register Read/Write
assign rvfi_rs1_addr  = rs1_addr_wb;
assign rvfi_rs1_rdata = rs1_rdata_wb;
assign rvfi_rs2_addr  = rs2_addr_wb;
assign rvfi_rs2_rdata = rs2_rdata_wb;
assign rvfi_rd_addr  = ((rd_dst_bank_wb == X_REG) && reg_wen_wb) ? (rd_addr_wb) : ('0);
assign rvfi_rd_wdata = (!rvfi_rd_addr) ? ('0) : (reg_wdata_wb);

// Program Counter
assign rvfi_pc_rdata = pc_wb;
assign rvfi_pc_wdata = pc_n_wb;

// Memory Access
assign rvfi_mem_addr  = mem_addr_wb;
assign rvfi_mem_rmask = mem_rmask_wb;
assign rvfi_mem_rdata = mem_rdata_wb;
assign rvfi_mem_wmask = mem_wmask_wb;
assign rvfi_mem_wdata = mem_wdata_wb;

// misa CSR
// wire [31:0] csr_mask_wb = {32{rvfi_valid_wb}};
wire [31:0] csr_rmask_wb = {32{rvfi_valid_wb}};
wire [31:0] csr_wmask_wb = {32{csr_wen_wb}};
assign rvfi_csr_misa_rmask = '1;
assign rvfi_csr_misa_rdata = misa;
assign rvfi_csr_misa_wmask = csr_wmask_wb;
assign rvfi_csr_misa_wdata = csr_wdata_wb;

`define assign_rvfi_csr(name) \
assign rvfi_csr_``name``_rmask = csr_rmask_wb; \
assign rvfi_csr_``name``_rdata = csr_rdata_wb; \
assign rvfi_csr_``name``_wmask = csr_wmask_wb; \
assign rvfi_csr_``name``_wdata = csr_wdata_wb;

`assign_rvfi_csr(mhartid)
`assign_rvfi_csr(mvendorid)
`assign_rvfi_csr(marchid)
`assign_rvfi_csr(mimpid)

`assign_rvfi_csr(mstatus)
`assign_rvfi_csr(mie)
`assign_rvfi_csr(mtvec)

`assign_rvfi_csr(mepc)
`assign_rvfi_csr(mcause)
`assign_rvfi_csr(mscratch)

`assign_rvfi_csr(fcsr)
`assign_rvfi_csr(fflags)
`assign_rvfi_csr(frm)


`default_nettype wire

endmodule
