///////////////////////////////////////////////////////////////////////////////////////////////////
//
//        CLASS: ls
//  DESCRIPTION: 
//         BUGS: ---
//       AUTHOR: Valmir F. Silva (), valmir.silva@ee.ufcg.edu.br
// ORGANIZATION: 
//      VERSION: 1.0
//      CREATED: 07/29/2024 07:37:29 PM
//     REVISION: ---
///////////////////////////////////////////////////////////////////////////////////////////////////
module mult(

            input logic         clock   ,
            input logic         nreset  ,
            input logic         valid   ,
            input logic [31:0]  a       ,
            input logic [31:0]  b       ,
            output logic [31:0] c       ,
            output logic ready          ,


  );

endmodule
