    
typedef enum bit {
    BAD_UVC_COV_ENABLE , 
    BAD_UVC_COV_DISABLE
} bad_uvc_cov_enable_enum;

typedef enum int {
    BAD_UVC_RST_STATE_PRE_RESET ,
    BAD_UVC_RST_STATE_IN_RESET  ,
    BAD_UVC_RST_STATE_POST_RESET
} bad_uvc_reset_state_enum;
