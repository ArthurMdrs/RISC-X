module OBI_controler #(
    parameter WIDTH = 32
) (
    OBI_if.MANAGER master
);
    

    


endmodule